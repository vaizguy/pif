
module pifctl (

    input  xclk   ,

    input  XI     ,
    output XO     ,
    
    output MiscReg
);

endmodule
