
module pifwb (

    inout  i2c_SCL,
    inout  i2c_SDA,

    input  xclk   ,

    output XI     ,
    input  XO
);

endmodule
